library verilog;
use verilog.vl_types.all;
entity genFace_vlg_check_tst is
    port(
        col_s0          : in     vl_logic;
        col_s1          : in     vl_logic;
        col_s2          : in     vl_logic;
        col_s3          : in     vl_logic;
        col_s4          : in     vl_logic;
        col_s5          : in     vl_logic;
        col_s6          : in     vl_logic;
        col_s7          : in     vl_logic;
        row_s0          : in     vl_logic;
        row_s1          : in     vl_logic;
        row_s2          : in     vl_logic;
        row_s3          : in     vl_logic;
        row_s4          : in     vl_logic;
        row_s5          : in     vl_logic;
        row_s6          : in     vl_logic;
        row_s7          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end genFace_vlg_check_tst;
