library verilog;
use verilog.vl_types.all;
entity CompareNum_vlg_vec_tst is
end CompareNum_vlg_vec_tst;
