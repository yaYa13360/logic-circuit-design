library verilog;
use verilog.vl_types.all;
entity createNum2_vlg_vec_tst is
end createNum2_vlg_vec_tst;
