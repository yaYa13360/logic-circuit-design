library verilog;
use verilog.vl_types.all;
entity projectFull_vlg_check_tst is
    port(
        gamest          : in     vl_logic;
        id0             : in     vl_logic;
        id1             : in     vl_logic;
        id2             : in     vl_logic;
        id3             : in     vl_logic;
        it0             : in     vl_logic;
        it1             : in     vl_logic;
        it2             : in     vl_logic;
        it3             : in     vl_logic;
        L1              : in     vl_logic;
        L2              : in     vl_logic;
        L3              : in     vl_logic;
        L4              : in     vl_logic;
        md0             : in     vl_logic;
        md1             : in     vl_logic;
        md2             : in     vl_logic;
        md3             : in     vl_logic;
        mt0             : in     vl_logic;
        mt1             : in     vl_logic;
        mt2             : in     vl_logic;
        mt3             : in     vl_logic;
        TFS1            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end projectFull_vlg_check_tst;
