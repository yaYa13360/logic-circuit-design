library verilog;
use verilog.vl_types.all;
entity projectFull_vlg_vec_tst is
end projectFull_vlg_vec_tst;
