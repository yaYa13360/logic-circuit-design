library verilog;
use verilog.vl_types.all;
entity projectFull_vlg_sample_tst is
    port(
        enter           : in     vl_logic;
        in0             : in     vl_logic;
        in1             : in     vl_logic;
        in2             : in     vl_logic;
        in3             : in     vl_logic;
        in4             : in     vl_logic;
        in5             : in     vl_logic;
        in6             : in     vl_logic;
        in7             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end projectFull_vlg_sample_tst;
