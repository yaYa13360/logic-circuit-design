library verilog;
use verilog.vl_types.all;
entity createNum2_vlg_sample_tst is
    port(
        clk1            : in     vl_logic;
        clk2            : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end createNum2_vlg_sample_tst;
