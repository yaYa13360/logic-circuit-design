library verilog;
use verilog.vl_types.all;
entity creatNum_vlg_vec_tst is
end creatNum_vlg_vec_tst;
