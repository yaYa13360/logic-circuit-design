library verilog;
use verilog.vl_types.all;
entity projectFull_vlg_sample_tst is
    port(
        enter           : in     vl_logic;
        g0              : in     vl_logic;
        g1              : in     vl_logic;
        g2              : in     vl_logic;
        g3              : in     vl_logic;
        g4              : in     vl_logic;
        g5              : in     vl_logic;
        g6              : in     vl_logic;
        g7              : in     vl_logic;
        mad0            : in     vl_logic;
        mad1            : in     vl_logic;
        mad2            : in     vl_logic;
        mad3            : in     vl_logic;
        mat0            : in     vl_logic;
        mat1            : in     vl_logic;
        mat2            : in     vl_logic;
        mat3            : in     vl_logic;
        mid0            : in     vl_logic;
        mid1            : in     vl_logic;
        mid2            : in     vl_logic;
        mid3            : in     vl_logic;
        mit0            : in     vl_logic;
        mit1            : in     vl_logic;
        mit2            : in     vl_logic;
        mit3            : in     vl_logic;
        restart         : in     vl_logic;
        start           : in     vl_logic;
        u0              : in     vl_logic;
        u1              : in     vl_logic;
        u2              : in     vl_logic;
        u3              : in     vl_logic;
        u4              : in     vl_logic;
        u5              : in     vl_logic;
        u6              : in     vl_logic;
        u7              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end projectFull_vlg_sample_tst;
