library verilog;
use verilog.vl_types.all;
entity creatNum_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        clk2            : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end creatNum_vlg_sample_tst;
