library verilog;
use verilog.vl_types.all;
entity genFace_vlg_vec_tst is
end genFace_vlg_vec_tst;
