library verilog;
use verilog.vl_types.all;
entity countLife_vlg_vec_tst is
end countLife_vlg_vec_tst;
