library verilog;
use verilog.vl_types.all;
entity projectFull is
    port(
        TFS0            : out    vl_logic;
        enter           : in     vl_logic;
        g0              : in     vl_logic;
        g1              : in     vl_logic;
        g2              : in     vl_logic;
        g3              : in     vl_logic;
        g4              : in     vl_logic;
        g5              : in     vl_logic;
        g6              : in     vl_logic;
        g7              : in     vl_logic;
        u0              : in     vl_logic;
        u1              : in     vl_logic;
        u2              : in     vl_logic;
        u3              : in     vl_logic;
        u4              : in     vl_logic;
        u5              : in     vl_logic;
        u6              : in     vl_logic;
        u7              : in     vl_logic;
        TFS1            : out    vl_logic
    );
end projectFull;
