library verilog;
use verilog.vl_types.all;
entity matrixFace_vlg_vec_tst is
end matrixFace_vlg_vec_tst;
