library verilog;
use verilog.vl_types.all;
entity projectFull_vlg_check_tst is
    port(
        TFS0            : in     vl_logic;
        TFS1            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end projectFull_vlg_check_tst;
